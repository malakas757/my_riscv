`timescale 1ns/1ps
import common::*;

module int1_alu_bju(/*AUTOARG*/
   // Outputs
   writeback2_valid, writeback2_need_to_wb, writeback2_prd,
   writeback2_robid, writeback2_data, ex2if_branch_valid,
   ex2if_branch_taken, ex2if_branch_addr, ex2if_branch_target_addr,
   ex2if_branch_update_GHSR, ex2if_GHSR_restore, branch_target_pc,
   branch_flush, branch_flush_robid,
   // Inputs
   clk, reset_n, flush_valid, flush_robid, int1_valid, int1_pc,
   int1_control, int1_rs1, int1_rs2, int1_T, int1_robid
   );
   input                       clk;
   input                       reset_n;
   input                       flush_valid;
   input [ROB_WIDTH:0] 	       flush_robid;

   //from buffer
   input                       int1_valid;
   input logic [31:0] 	       int1_pc;
   input control_type          int1_control;
   input logic [31:0]          int1_rs1;
   input logic [31:0]          int1_rs2;
   input logic [PRF_WIDTH-1:0] int1_T;
   input logic [ROB_WIDTH:0]   int1_robid;
   //output to writeback2 alu
   output logic                 writeback2_valid;//int0 mul
   output logic 		writeback2_need_to_wb;
   output logic [PRF_WIDTH-1:0] writeback2_prd;                     
   output logic [ROB_WIDTH:0] 	writeback2_robid;                     
   output logic [31:0] 		writeback2_data;  

   //output about bp
   output  logic 		            ex2if_branch_valid;   // remeber comb with valid
   output  logic 			    ex2if_branch_taken;
   output  logic [31:0] 		    ex2if_branch_addr;//pc
   output  logic [31:0] 		    ex2if_branch_target_addr;//branch target pc,this used to update btb  
   output  logic 			    ex2if_branch_update_GHSR; //
   output  logic [GSHARE_GHSR_WIDTH-1:0]    ex2if_GHSR_restore ;
   output  logic [31:0] 		    branch_target_pc; // branch target pc(after latch),this is used to redirect
   output  logic 			    branch_flush;//after latch ,need to input back to this module   
   output  logic [ROB_WIDTH:0] 		    branch_flush_robid;//after latch ,need to input back to this module   



   logic [31:0] 		alu_left_operand;
   logic [31:0] 		alu_right_operand;


   logic                        is_bj;
   
   //these are results generated by bju
   logic                        bju_flush_result;// is just cal result need comb with valid
   logic                        bju_branch_taken;//
   logic                        bju_branch_update_GHSR;//
   logic [31:0] 		bju_branch_target_pc;//
   logic [GSHARE_GHSR_WIDTH-1:0]    bju_GHSR_restore ;
   logic [31:0] 		j_next_pc;// result for jal and jalr next pc
   logic [31:0] 		alu_data;// result for alu_data

   //wb reg
   logic 			wb_reg_valid;
   logic 			wb_reg_need_to_wb;
   logic [PRF_WIDTH-1:0] 	wb_reg_prd;                     
   logic [ROB_WIDTH:0] 		wb_reg_robid;                     
   logic [31:0] 		wb_reg_data;
   logic 			wb_need_to_flush;

   
   //latch the flush information
  // logic                        branch_flush_latch;
  // logic                        branch_taken_latch;
  // logic                        branch_valid_latch;
  // logic [31:0] 		branch_target_pc_latch;
  // logic [ROB_WIDTH:0] 		branch_flush_robid_latch;
  // logic [31:0] 		branch_pc_latch;//used to update btb
  // logic 			branch_update_GHSR_latch; //
  // logic [GSHARE_GHSR_WIDTH-1:0] GHSR_restore_latch ;
   


   assign is_bj = int1_control.is_jump | int1_control.is_jumpr | int1_control.is_branch;


   

   always_comb begin: operand_selector
      alu_left_operand  = (int1_control.is_auipc)? int1_pc : int1_rs1 ;// add AUIPC
      alu_right_operand = int1_rs2;
      if (int1_control.alu_src) begin
         alu_right_operand = int1_control.imm_data;
      end
   end



   
   //for alu
   alu inst_alu(
		.control(int1_control.alu_op),
		.left_operand(alu_left_operand), 
		.right_operand(alu_right_operand),
		.result(alu_data)
		);


   


   //bju


        //latch the flush infor
        always_ff@(posedge clk) begin
	   if (~reset_n | flush_valid) begin
	      branch_flush      <= '0; 
	      branch_flush_robid      <= '0; 
	    //  branch_taken_latch      = '0; 
	    //  branch_valid_latch      = '0; 
	      branch_target_pc  <= '0;  	      
	   //   branch_pc_latch  = '0;  	      
	   //   branch_update_GHSR_latch       = '0; 	      
	   //   GHSR_restore_latch       = '0; 	      
	   end
	   else begin
	      branch_flush            <= int1_valid & bju_flush_result; 
	      branch_flush_robid      <= int1_robid; 
	   //   branch_taken_latch      = bju_branch_taken; 
	   //  branch_valid_latch      = int1_valid & is_bj; 
	      branch_target_pc        <= bju_branch_target_pc;  	      
	   //   branch_pc_latch         = int1_pc;  	      
	   //   branch_update_GHSR_latch = int1_valid & bju_branch_update_GHSR; 	     
	   //   GHSR_restore_latch       = bju_GHSR_restore; 	      
	   end // else: !if(~reset_n & need_to_flush)
	end


   
   bju inst_bju(
		// Outputs
		.j_next_pc		(j_next_pc[31:0]),
		.branch_target_pc	(bju_branch_target_pc),
		.branch_taken		(bju_branch_taken),
		.flush			(bju_flush_result),
		.GHSR_restore		(bju_GHSR_restore),
		.update_GHSR		(bju_branch_update_GHSR),
		// Inputs
		.left_operand		(int1_rs1),
		.right_operand		(int1_rs2),
		.pc			(int1_pc),
		.clk			(clk),
		.reset_n		(reset_n),
		.control		(int1_control),
		.immediate_data		(int1_control.imm_data),
		.branch_predict		(int1_control.predict));


   assign  ex2if_branch_addr        = int1_pc;
   assign  ex2if_branch_valid       = int1_valid & is_bj & ~flush_valid;   // remeber comb with valid
   assign  ex2if_branch_taken       = bju_branch_taken; 
   assign  ex2if_branch_target_addr = bju_branch_target_pc; // branch target pc,this used to update btb
   assign  ex2if_branch_update_GHSR = int1_valid & bju_branch_update_GHSR & ~flush_valid; //
   assign  ex2if_GHSR_restore       = bju_GHSR_restore;
 //  assign  branch_target_pc         = branch_target_pc_latch; // branch target pc
 //  assign  branch_flush             = branch_flush_latch;     


   //wb
   assign wb_need_to_flush = (flush_valid & (wb_reg_robid[ROB_WIDTH] ^ flush_robid[ROB_WIDTH] ^ (wb_reg_robid[ROB_WIDTH-1:0] > flush_robid[ROB_WIDTH-1:0])))?1:0;
   assign writeback2_need_to_wb  = wb_reg_need_to_wb;
   assign writeback2_valid       = wb_reg_valid & ~flush_valid;
   assign writeback2_prd         = wb_reg_prd;
   assign writeback2_robid       = wb_reg_robid;
   assign writeback2_data        = wb_reg_data;
   
   
   always_ff@(posedge clk) begin
      if(~reset_n | wb_need_to_flush) begin
	 wb_reg_valid      <= 1'b0;
	 wb_reg_robid      <= '0;
	 wb_reg_prd        <= '0;
	 wb_reg_data       <= '0;
	 wb_reg_need_to_wb <= '0;
      end
      else if ( ~flush_valid ) begin
	 wb_reg_valid      <= int1_valid;
	 wb_reg_robid      <= int1_robid;
	 wb_reg_prd        <= int1_T;
	 wb_reg_data       <= (int1_control.is_jumpr | int1_control.is_jump)? j_next_pc : alu_data;
	 wb_reg_need_to_wb <= int1_control.reg_write;	 
      end	 
   end
   
endmodule
