`timescale 1ns / 1ps

import common::*;


module test(
/*AUTOARG*/
   // Outputs
   out,
   // Inputs
   in
   );
   input in;

   output out;
   
endmodule
