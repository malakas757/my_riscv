package common;


   

   
endpackage
