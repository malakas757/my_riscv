`timescale 1ns/1ps

import common::*;

module int0_alu_mul(/*AUTOARG*/);
   

   







   

endmodule // int0_alu_mul
