`timescale 1ns/1ps
import common::*;

module int0_mul_alu(/*AUTOARG*/
   // Outputs
   mul_is_busy, writeback0_valid, writeback0_need_to_wb,
   writeback0_prd, writeback0_robid, writeback0_data,
   writeback1_valid, writeback1_need_to_wb, writeback1_robid,
   writeback1_prd, writeback1_data,
   // Inputs
   clk, reset_n, flush_valid, flush_robid, int0_valid, int0_pc,
   int0_control, int0_rs1, int0_rs2, int0_T, int0_robid
   );

   input                       clk;
   input                       reset_n;
   input                       flush_valid;
   input [ROB_WIDTH:0] 	       flush_robid;
   output 		       mul_is_busy;//always 1 because pipeline mul unit
   
   

   input                       int0_valid;
   input logic [31:0] 	       int0_pc;
   input control_type          int0_control;
   input logic [31:0]          int0_rs1;
   input logic [31:0]          int0_rs2;
   input logic [PRF_WIDTH-1:0] int0_T;
   input logic [ROB_WIDTH:0]   int0_robid;


   //output to mul_wb
   output logic                 writeback0_valid;//int0 mul
   output logic 		writeback0_need_to_wb;
   output logic [PRF_WIDTH-1:0] writeback0_prd;                     
   output logic [ROB_WIDTH:0] 	writeback0_robid;                     
   output logic [31:0] 		writeback0_data;                     
   //output to alu_wb
   output logic                 writeback1_valid;//int0 mul
   output logic 		writeback1_need_to_wb;
   output logic [ROB_WIDTH:0] 	writeback1_robid;
   output logic [PRF_WIDTH-1:0] writeback1_prd;                     
   output logic [31:0] 		writeback1_data;


   logic [31:0] 		left_operand;
   logic [31:0] 		right_operand;
   logic [63:0] 		mul_out_data;
   logic 			mul_done;
   logic 			mul_out_valid;
   logic [ROB_WIDTH:0] 		mul_out_robid;
   logic [PRF_WIDTH-1:0] 	mul_out_T;

   



   
   always_comb begin: operand_selector
      left_operand  = (int0_control.is_auipc)? int0_pc : int0_rs1 ;// add AUIPC
      right_operand = int0_rs2;
      if (int0_control.alu_src) begin
         right_operand = int0_control.imm_data;
      end
   end

   //for alu
   alu inst_alu(
		.control(int0_control.alu_op),
		.left_operand(left_operand), 
		.right_operand(right_operand),
		.result(writeback1_data)
		);

   assign writeback1_need_to_wb = int0_control.reg_write;
   assign writeback1_valid =  ~flush_valid & int0_valid & ~int0_control.is_mul;
   assign writeback1_prd = int0_T;
   assign writeback1_robid = int0_robid;

   //for mul
   mult inst_mult(
		  // Outputs
		  .product		(mul_out_data),
		  .done			(mul_done),
		  .out_valid		(mul_out_valid),
		  .out_rob_id		(mul_out_robid),
		  .out_prf_id		(mul_out_T),
		  // Inputs
		  .clock		(clk),
		  .reset		(~reset_n),
		  .start		(int0_control.is_mul & int0_valid),
		  .sign			(2'b11),// only support MUL,so should be signed
		  .mcand		(left_operand),
		  .mplier		(right_operand),
		  .valid		(int0_control.is_mul & int0_valid),
		  .rob_id		(int0_robid),
		  .flush_robid		(flush_robid[ROB_WIDTH:0]),
		  .prf_id		(int0_T),
		  .flush_valid		(flush_valid));
   
   assign writeback0_data = mul_out_data[31:0];
   assign writeback0_valid = mul_done & mul_out_valid;
   assign writeback0_prd = mul_out_T;
   assign writeback0_robid = mul_out_robid;
   assign writeback0_need_to_wb = 1'b1;//mul must be a reg write instr
   assign mul_is_busy = 1'b0;
  
   


endmodule

