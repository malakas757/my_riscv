//system
`define   ADDR_WIDTH        32
//cache  
`define   CACHELINE_WIDTH   512  
`define   CACHE_SET         64
`define   CACHE_TAG_WIDTH   20 // 32-log(512/8)-log(64)
//
`define   INSTR_WIDTH       8 // 32-log(512/8)-log(64)      

