`define ROB_WIDTH   7 // 2 bits(3 chn) + 2bits(4 banks) + 3bits(SWB_DEPTH)
`define ROB_WIDTH   7 // 2 bits(3 chn) + 2bits(4 banks) + 3bits(SWB_DEPTH)
