`timescale 1ns/1ps

import common::*;


module int2_lsu(/*AUTOARG*/);

   








endmodule
